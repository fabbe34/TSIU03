library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; 
use work.common.all;

library work;

entity TB_equ is


end entity;

Architecture sim of TB_equ is

-- dut signals
	signal clk,rstn : std_logic:='1';
	signal x_in : signed(15 downto 0) := "0101010101010101";
	signal coeff : coefficients:=
 (X"0003", -- mem(A0) = 5,52345897316551E-05
  X"0004", -- mem(A1) = 6,80644238118407E-05
  X"0005", -- mem(A2) = 8,24589475370423E-05
  X"0006", -- mem(A3) = 9,84452601078052E-05
  X"0007", -- mem(A4) = 0,000116068950190736
  X"0008", -- mem(A5) = 0,000135248483153016
  X"000A", -- mem(A6) = 0,000155968483382642
  X"000B", -- mem(A7) = 0,000178155643529953
  X"000D", -- mem(A8) = 0,000201821969265627
  X"000E", -- mem(A9) = 0,000226791245218498
  X"0010", -- mem(A10) = 0,000252911486259129
  X"0012", -- mem(A11) = 0,000279962554194093
  X"0014", -- mem(A12) = 0,00030793593714325
  X"0016", -- mem(A13) = 0,000336384341656877
  X"0017", -- mem(A14) = 0,00036505315389209
  X"0019", -- mem(A15) = 0,000393764380603094
  X"001B", -- mem(A16) = 0,000421962671475817
  X"001D", -- mem(A17) = 0,000449453667631933
  X"001F", -- mem(A18) = 0,00047571587913539
  X"0020", -- mem(A19) = 0,000500356402770411
  X"0022", -- mem(A20) = 0,000522832192503619
  X"0023", -- mem(A21) = 0,000542673488164318
  X"0024", -- mem(A22) = 0,000559329327434486
  X"0025", -- mem(A23) = 0,000572241709785608
  X"0026", -- mem(A24) = 0,000580814114668601
  X"0026", -- mem(A25) = 0,000584487717924256
  X"0026", -- mem(A26) = 0,00058265572366315
  X"0025", -- mem(A27) = 0,000574688639465408
  X"0024", -- mem(A28) = 0,000560044620486117
  X"0023", -- mem(A29) = 0,000538073861900304
  X"0021", -- mem(A30) = 0,00050821343574349
  X"001E", -- mem(A31) = 0,000469925491451767
  X"001B", -- mem(A32) = 0,000422660047205058
  X"0018", -- mem(A33) = 0,000365954198445497
  X"0013", -- mem(A34) = 0,000299335869329561
  X"000E", -- mem(A35) = 0,000222443384258505
  X"0008", -- mem(A36) = 0,000134921514874078
  X"0002", -- mem(A37) = 3,65225417273913E-05
  X"FFFB", -- mem(A38) = -7,29493426174901E-05
  X"FFF3", -- mem(A39) = -0,000193587399621588
  X"FFEA", -- mem(A40) = -0,000325432202961925
  X"FFE1", -- mem(A41) = -0,00046837665772445
  X"FFD7", -- mem(A42) = -0,000622245244910659
  X"FFCC", -- mem(A43) = -0,000786758526926491
  X"FFC1", -- mem(A44) = -0,000961489229025817
  X"FFB4", -- mem(A45) = -0,00114593048250338
  X"FFA8", -- mem(A46) = -0,00133942150087028
  X"FF9B", -- mem(A47) = -0,00154119322655691
  X"FF8D", -- mem(A48) = -0,00175034293294687
  X"FF7F", -- mem(A49) = -0,00196584098315754
  X"FF70", -- mem(A50) = -0,00218654338994281
  X"FF62", -- mem(A51) = -0,00241115761968007
  X"FF53", -- mem(A52) = -0,00263828709212596
  X"FF44", -- mem(A53) = -0,00286640623694068
  X"FF35", -- mem(A54) = -0,00309388163147455
  X"FF26", -- mem(A55) = -0,00331895035035988
  X"FF18", -- mem(A56) = -0,00353977941381046
  X"FF0A", -- mem(A57) = -0,00375440536325517
  X"FEFC", -- mem(A58) = -0,00396080625689552
  X"FEEF", -- mem(A59) = -0,00415687914875703
  X"FEE3", -- mem(A60) = -0,00434045401858865
  X"FED8", -- mem(A61) = -0,00450932118459746
  X"FECE", -- mem(A62) = -0,004661223153316
  X"FEC5", -- mem(A63) = -0,00479389935618745
  X"FEBE", -- mem(A64) = -0,00490507014977938
  X"FEB8", -- mem(A65) = -0,00499247327398246
  X"FEB4", -- mem(A66) = -0,00505387509139222
  X"FEB2", -- mem(A67) = -0,00508708333639423
  X"FEB2", -- mem(A68) = -0,0050899675300111
  X"FEB4", -- mem(A69) = -0,00506048149787073
  X"FEB8", -- mem(A70) = -0,00499667755645861
  X"FEBF", -- mem(A71) = -0,00489671178382397
  X"FEC8", -- mem(A72) = -0,00475889570663942
  X"FED3", -- mem(A73) = -0,00458167039531877
  X"FEE2", -- mem(A74) = -0,0043636636512899
  X"FEF3", -- mem(A75) = -0,00410367271627798
  X"FF06", -- mem(A76) = -0,0038007026511583
  X"FF1D", -- mem(A77) = -0,00345396875335889
  X"FF37", -- mem(A78) = -0,00306290894816429
  X"FF53", -- mem(A79) = -0,002627208017236
  X"FF73", -- mem(A80) = -0,00214679032613268
  X"FF95", -- mem(A81) = -0,0016218413607925
  X"FFBB", -- mem(A82) = -0,00105280860114309
  X"FFE3", -- mem(A83) = -0,000440415747913956
  X"000E", -- mem(A84) = 0,000214348841593246
  X"003B", -- mem(A85) = 0,000910212246140831
  X"006B", -- mem(A86) = 0,00164562954448378
  X"009E", -- mem(A87) = 0,00241878466850675
  X"00D3", -- mem(A88) = 0,00322758294957264
  X"010A", -- mem(A89) = 0,00406967719689579
  X"0143", -- mem(A90) = 0,00494245190402161
  X"017E", -- mem(A91) = 0,00584306053996237
  X"01BB", -- mem(A92) = 0,00676841032562725
  X"01F9", -- mem(A93) = 0,0077151960908742
  X"0238", -- mem(A94) = 0,00867990633312393
  X"0279", -- mem(A95) = 0,00965884386650041
  X"02B9", -- mem(A96) = 0,0106481450039346
  X"02FB", -- mem(A97) = 0,0116437993071172
  X"033C", -- mem(A98) = 0,0126416752627509
  X"037D", -- mem(A99) = 0,0136375336043661
  X"03BE", -- mem(A100) = 0,0146270693199103
  X"03FE", -- mem(A101) = 0,0156059169605172
  X"043D", -- mem(A102) = 0,0165696934074244
  X"047B", -- mem(A103) = 0,0175140124354336
  X"04B8", -- mem(A104) = 0,0184345177588436
  X"04F2", -- mem(A105) = 0,0193269121662617
  X"052B", -- mem(A106) = 0,0201869747913066
  X"0561", -- mem(A107) = 0,0210106033949866
  X"0594", -- mem(A108) = 0,021793822063175
  X"05C4", -- mem(A109) = 0,0225328251194889
  X"05F2", -- mem(A110) = 0,0232239869415944
  X"061B", -- mem(A111) = 0,0238638992862979
  X"0642", -- mem(A112) = 0,0244493809839418
  X"0664", -- mem(A113) = 0,0249775077650079
  X"0683", -- mem(A114) = 0,0254456290995872
  X"069E", -- mem(A115) = 0,025851381584397
  X"06B4", -- mem(A116) = 0,0261927156120729
  X"06C6", -- mem(A117) = 0,026467893094339
  X"06D4", -- mem(A118) = 0,026675516869461
  X"06DD", -- mem(A119) = 0,0268145235502832
  X"06E1", -- mem(A120) = 0,0268842055657813
  X"06E1", -- mem(A121) = 0,0268842055657813
  X"06DD", -- mem(A122) = 0,0268145235502832
  X"06D4", -- mem(A123) = 0,026675516869461
  X"06C6", -- mem(A124) = 0,026467893094339
  X"06B4", -- mem(A125) = 0,0261927156120729
  X"069E", -- mem(A126) = 0,025851381584397
  X"0683", -- mem(A127) = 0,0254456290995872
  X"0664", -- mem(A128) = 0,0249775077650079
  X"0642", -- mem(A129) = 0,0244493809839418
  X"061B", -- mem(A130) = 0,0238638992862979
  X"05F2", -- mem(A131) = 0,0232239869415944
  X"05C4", -- mem(A132) = 0,0225328251194889
  X"0594", -- mem(A133) = 0,021793822063175
  X"0561", -- mem(A134) = 0,0210106033949866
  X"052B", -- mem(A135) = 0,0201869747913066
  X"04F2", -- mem(A136) = 0,0193269121662617
  X"04B8", -- mem(A137) = 0,0184345177588436
  X"047B", -- mem(A138) = 0,0175140124354336
  X"043D", -- mem(A139) = 0,0165696934074244
  X"03FE", -- mem(A140) = 0,0156059169605172
  X"03BE", -- mem(A141) = 0,0146270693199103
  X"037D", -- mem(A142) = 0,0136375336043661
  X"033C", -- mem(A143) = 0,0126416752627509
  X"02FB", -- mem(A144) = 0,0116437993071172
  X"02B9", -- mem(A145) = 0,0106481450039346
  X"0279", -- mem(A146) = 0,00965884386650041
  X"0238", -- mem(A147) = 0,00867990633312393
  X"01F9", -- mem(A148) = 0,0077151960908742
  X"01BB", -- mem(A149) = 0,00676841032562725
  X"017E", -- mem(A150) = 0,00584306053996237
  X"0143", -- mem(A151) = 0,00494245190402161
  X"010A", -- mem(A152) = 0,00406967719689579
  X"00D3", -- mem(A153) = 0,00322758294957264
  X"009E", -- mem(A154) = 0,00241878466850675
  X"006B", -- mem(A155) = 0,00164562954448378
  X"003B", -- mem(A156) = 0,000910212246140831
  X"000E", -- mem(A157) = 0,000214348841593246
  X"FFE3", -- mem(A158) = -0,000440415747913956
  X"FFBB", -- mem(A159) = -0,00105280860114309
  X"FF95", -- mem(A160) = -0,0016218413607925
  X"FF73", -- mem(A161) = -0,00214679032613268
  X"FF53", -- mem(A162) = -0,002627208017236
  X"FF37", -- mem(A163) = -0,00306290894816429
  X"FF1D", -- mem(A164) = -0,00345396875335889
  X"FF06", -- mem(A165) = -0,0038007026511583
  X"FEF3", -- mem(A166) = -0,00410367271627798
  X"FEE2", -- mem(A167) = -0,0043636636512899
  X"FED3", -- mem(A168) = -0,00458167039531877
  X"FEC8", -- mem(A169) = -0,00475889570663942
  X"FEBF", -- mem(A170) = -0,00489671178382397
  X"FEB8", -- mem(A171) = -0,00499667755645861
  X"FEB4", -- mem(A172) = -0,00506048149787073
  X"FEB2", -- mem(A173) = -0,0050899675300111
  X"FEB2", -- mem(A174) = -0,00508708333639423
  X"FEB4", -- mem(A175) = -0,00505387509139222
  X"FEB8", -- mem(A176) = -0,00499247327398246
  X"FEBE", -- mem(A177) = -0,00490507014977938
  X"FEC5", -- mem(A178) = -0,00479389935618745
  X"FECE", -- mem(A179) = -0,004661223153316
  X"FED8", -- mem(A180) = -0,00450932118459746
  X"FEE3", -- mem(A181) = -0,00434045401858865
  X"FEEF", -- mem(A182) = -0,00415687914875703
  X"FEFC", -- mem(A183) = -0,00396080625689552
  X"FF0A", -- mem(A184) = -0,00375440536325517
  X"FF18", -- mem(A185) = -0,00353977941381046
  X"FF26", -- mem(A186) = -0,00331895035035988
  X"FF35", -- mem(A187) = -0,00309388163147455
  X"FF44", -- mem(A188) = -0,00286640623694068
  X"FF53", -- mem(A189) = -0,00263828709212596
  X"FF62", -- mem(A190) = -0,00241115761968007
  X"FF70", -- mem(A191) = -0,00218654338994281
  X"FF7F", -- mem(A192) = -0,00196584098315754
  X"FF8D", -- mem(A193) = -0,00175034293294687
  X"FF9B", -- mem(A194) = -0,00154119322655691
  X"FFA8", -- mem(A195) = -0,00133942150087028
  X"FFB4", -- mem(A196) = -0,00114593048250338
  X"FFC1", -- mem(A197) = -0,000961489229025817
  X"FFCC", -- mem(A198) = -0,000786758526926491
  X"FFD7", -- mem(A199) = -0,000622245244910659
  X"FFE1", -- mem(A200) = -0,00046837665772445
  X"FFEA", -- mem(A201) = -0,000325432202961925
  X"FFF3", -- mem(A202) = -0,000193587399621588
  X"FFFB", -- mem(A203) = -7,29493426174901E-05
  X"0002", -- mem(A204) = 3,65225417273913E-05
  X"0008", -- mem(A205) = 0,000134921514874078
  X"000E", -- mem(A206) = 0,000222443384258505
  X"0013", -- mem(A207) = 0,000299335869329561
  X"0018", -- mem(A208) = 0,000365954198445497
  X"001B", -- mem(A209) = 0,000422660047205058
  X"001E", -- mem(A210) = 0,000469925491451767
  X"0021", -- mem(A211) = 0,00050821343574349
  X"0023", -- mem(A212) = 0,000538073861900304
  X"0024", -- mem(A213) = 0,000560044620486117
  X"0025", -- mem(A214) = 0,000574688639465408
  X"0026", -- mem(A215) = 0,00058265572366315
  X"0026", -- mem(A216) = 0,000584487717924256
  X"0026", -- mem(A217) = 0,000580814114668601
  X"0025", -- mem(A218) = 0,000572241709785608
  X"0024", -- mem(A219) = 0,000559329327434486
  X"0023", -- mem(A220) = 0,000542673488164318
  X"0022", -- mem(A221) = 0,000522832192503619
  X"0020", -- mem(A222) = 0,000500356402770411
  X"001F", -- mem(A223) = 0,00047571587913539
  X"001D", -- mem(A224) = 0,000449453667631933
  X"001B", -- mem(A225) = 0,000421962671475817
  X"0019", -- mem(A226) = 0,000393764380603094
  X"0017", -- mem(A227) = 0,00036505315389209
  X"0016", -- mem(A228) = 0,000336384341656877
  X"0014", -- mem(A229) = 0,00030793593714325
  X"0012", -- mem(A230) = 0,000279962554194093
  X"0010", -- mem(A231) = 0,000252911486259129
  X"000E", -- mem(A232) = 0,000226791245218498
  X"000D", -- mem(A233) = 0,000201821969265627
  X"000B", -- mem(A234) = 0,000178155643529953
  X"000A", -- mem(A235) = 0,000155968483382642
  X"0008", -- mem(A236) = 0,000135248483153016
  X"0007", -- mem(A237) = 0,000116068950190736
  X"0006", -- mem(A238) = 9,84452601078052E-05
  X"0005", -- mem(A239) = 8,24589475370423E-05
  X"0004", -- mem(A240) = 6,80644238118407E-05
  X"0003", -- mem(A241) = 5,52345897316551E-05
  X"0007"); -- mem(A242) = 0,000113538734273173)
  
  
  signal done : boolean := false;
  
  
  
  component FIR_PE is
	port(
	
		clk, rstn : in std_logic;
			--start   	 : in std_logic;
			x_in 		 : in signed(15 downto 0);
			y_out		 : out signed(15 downto 0);
			coeff 	 : in coefficients
		);
	end component;
	
	
begin 


	clk <= not clk after 10ns when not done;
	rstn <= '0', '1' after 50 ns;
	done <= false, true after 1 ms;

	
	end architecture;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; 
use ieee.math_real.all;


package Common is

	type coefficients is array (0 to 255) of signed(15 downto 0);
	
	type input_memory is array (0 to 255) of signed (15 downto 0);
	
	end Common;
	
	
	
	package body Common is 
	
	
	end common;
	
	